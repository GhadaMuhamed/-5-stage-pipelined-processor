
LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

ENTITY mux2 IS  
Generic (n : integer :=16);
PORT (
IN1,IN2: IN STD_LOGIC_VECTOR(n-1 DOWNTO 0);
SEl:IN STD_LOGIC;
OUT1:OUT  STD_LOGIC_VECTOR(n-1 DOWNTO 0)
);    
END ENTITY mux2;


ARCHITECTURE ArchMux OF mux2 IS
BEGIN
OUT1 <= IN1 WHEN SEl='0'
ELSE IN2;
END ArchMux;